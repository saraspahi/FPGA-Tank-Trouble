/************************************************************************
Avalon-MM Interface VGA Text mode display

Register Map:
0x000-0x0257 : VRAM, 80x30 (2400 byte, 600 word) raster order (first column then row)
0x258        : control register

VRAM Format:
X->
[ 31  30-24][ 23  22-16][ 15  14-8 ][ 7    6-0 ]
[IV3][CODE3][IV2][CODE2][IV1][CODE1][IV0][CODE0]

IVn = Draw inverse glyph
CODEn = Glyph code from IBM codepage 437

Control Register Format:
[[31-25][24-21][20-17][16-13][ 12-9][ 8-5 ][ 4-1 ][   0    ] 
[[RSVD ][FGD_R][FGD_G][FGD_B][BKG_R][BKG_G][BKG_B][RESERVED]

VSYNC signal = bit which flips on every Vsync (time for new frame), used to synchronize software
BKG_R/G/B = Background color, flipped with foreground when IVn bit is set
FGD_R/G/B = Foreground color, flipped with background when Inv bit is set

************************************************************************/
`define NUM_REGS 601 //80*30 characters / 4 characters per register
`define CTRL_REG 600 //index of control register

module vga_text_avl_interface (
	// Avalon Clock Input, note this clock is also used for VGA, so this must be 50Mhz
	// We can put a clock divider here in the future to make this IP more generalizable
	input logic CLK,
	
	// Avalon Reset Input
	input logic RESET,
	
	// Avalon-MM Slave Signals
	input  logic AVL_READ,					// Avalon-MM Read
	input  logic AVL_WRITE,					// Avalon-MM Write
	input  logic AVL_CS,					// Avalon-MM Chip Select
	input  logic [3:0] AVL_BYTE_EN,			// Avalon-MM Byte Enable
	input  logic [11:0] AVL_ADDR,			// Avalon-MM Address
	input  logic [31:0] AVL_WRITEDATA,		// Avalon-MM Write Data
	output logic [31:0] AVL_READDATA,		// Avalon-MM Read Data
	
	// Exported Conduit (mapped to VGA port - make sure you export in Platform Designer)
	output logic [3:0]  red, green, blue,	// VGA color channels (mapped to output pins in top-level)
	output logic hs, vs						// VGA HS/VS
);

logic [31:0] COLOR_REGS [8]; // Registers
//// Read and write from AVL interface to register block, note that READ waitstate = 1, so this should be in always_ff
//// implement control 
//always_comb
//begin
//	COLOR_REGS [0][31:0] = 32'h00000000;
//	COLOR_REGS [1][31:0] = 32'h00000014;
//	COLOR_REGS [2][31:0] = 32'hFFFFFF0F;
//	COLOR_REGS [3][31:0] = 32'hFF0F0FFF;
//	COLOR_REGS [4][31:0] = 32'hFFFF0FF0;
//	COLOR_REGS [5][31:0] = 32'hFFF0F0FF;
//	COLOR_REGS [6][31:0] = 32'hFF0FFFFF;
//	COLOR_REGS [7][31:0] = 32'hFF0FF0FF;
//end
//
always_ff@(posedge CLK)
begin 
if(AVL_WRITE && AVL_CS && AVL_ADDR[11])
begin

	COLOR_REGS[AVL_ADDR[2:0]][31:0] <= AVL_WRITEDATA[31:0];
	
end

if(AVL_READ && AVL_CS && AVL_ADDR[11])
begin
	//AVL_READDATA = COLOR_REGS[AVL_ADDR[2:0]];
end

else if(RESET)
	begin
		for(int i = 0; i<8; i++)
		begin
			//COLOR_REGS[i] <= 32'hFFFFFFF;
		end
	end
end
 
//put other local variables here
logic [31:0] Ram_Out;
logic [10:0] Font_Rom_ADDR;
logic [7:0]  Font_Rom_DATA;
logic [9:0]  DrawX, DrawY, Word_ADDR, Read_ADDR;
logic [11:0] Byte_ADDR;
logic [7:0] CodeN;
logic [31:0] LOCAL_REG, DATA_OUT;
logic [2:0] FONTR_I;
logic blank, PIX_CLK;
logic [3:0] FGD_I, BKG_I, FGD_R, FGD_B, FGD_G, BKG_R, BKG_B, BKG_G;

//logic [1:0] Byte_INDEX;
//logic CurrInv;
//Declare submodules..e.g. VGA controller, ROMS, etc

always_comb
begin
if(AVL_READ && AVL_CS)
	Read_ADDR = AVL_ADDR;
else
	Read_ADDR = Word_ADDR;
end

//always_comb
//
//begin
//if(AVL_ADDR[11])
//	AVL_READDATA = COLOR_REGS[AVL_ADDR[2:0]];
//else
//	AVL_READDATA = Ram_Out;
//end


ram1 ram1(.byteena_a(AVL_BYTE_EN), .clock(CLK), .data(AVL_WRITEDATA), .rdaddress(Read_ADDR),
			.wraddress(AVL_ADDR), .wren(AVL_WRITE && AVL_CS && ~AVL_ADDR[11]), .q(AVL_READDATA));

font_rom FR(.addr(Font_Rom_ADDR), .data(Font_Rom_DATA));
vga_controller VGA_C(.Clk(CLK), .Reset(RESET), .pixel_clk(PIX_CLK), .hs(hs), .vs(vs), .DrawX(DrawX), .DrawY(DrawY), .blank(blank)); 


// Give the Control Register Values
color_mapper CM(.DrawX(~DrawX[2:0]), .CLK(PIX_CLK), .Font_Rom_DATA(Font_Rom_DATA), .blank(blank),
						.FGD_R(FGD_R), .FGD_G(FGD_G), 
														.FGD_B(FGD_B), .BKG_R(BKG_R), 
														.BKG_G(BKG_G), .BKG_B(BKG_B),
														.INV(CodeN[7]), .Red(red), .Green(green), .Blue(blue)); 


														
//handle drawing (may either be combinational or sequential - or both).

	// Handle reading the Codes from the Local regs
always_comb
begin
	Byte_ADDR[11:0] = DrawX[9:3] + DrawY[9:4]*7'd80;
 	Word_ADDR = Byte_ADDR[11:1];
	
	if(Byte_ADDR[0] == 1'b0)
	begin
		CodeN[7:0] = AVL_READDATA[15:8];
		FGD_I[3:0] = AVL_READDATA[7:4];
		BKG_I[3:0] = AVL_READDATA[3:0];
	end
	
	else if(Byte_ADDR[0] == 1'b1)
	begin
		CodeN[7:0] = AVL_READDATA[31:24];
		FGD_I[3:0] = AVL_READDATA[23:20];
		BKG_I[3:0] = AVL_READDATA[19:16];		
	end
			
	else
	begin
		CodeN[7:0] = 8'h00;	
		FGD_I[3:0] = AVL_READDATA[23:20];
		BKG_I[3:0] = AVL_READDATA[19:16];
	end
	
	Font_Rom_ADDR = {{CodeN[6:0]}, {DrawY[3:0]}};
end

always_comb
begin
	if(FGD_I[0] == 1'b0)
	begin 
		FGD_R = COLOR_REGS[FGD_I[3:1]][12:9];
		FGD_G = COLOR_REGS[FGD_I[3:1]][8:5];
		FGD_B = COLOR_REGS[FGD_I[3:1]][4:1];
	end
	
	else
	begin 
		FGD_R = COLOR_REGS[FGD_I[3:1]][24:21];
		FGD_G = COLOR_REGS[FGD_I[3:1]][20:17];
		FGD_B = COLOR_REGS[FGD_I[3:1]][16:13];
	end
end

always_comb
begin
	if(BKG_I[0] == 1'b0)
	begin 
		BKG_R = COLOR_REGS[BKG_I[3:1]][12:9];
		BKG_G = COLOR_REGS[BKG_I[3:1]][8:5];
		BKG_B = COLOR_REGS[BKG_I[3:1]][4:1];
	end
	
	else
	begin 
		BKG_R = COLOR_REGS[BKG_I[3:1]][24:21];
		BKG_G = COLOR_REGS[BKG_I[3:1]][20:17];
		BKG_B = COLOR_REGS[BKG_I[3:1]][16:13];
	end
end

endmodule