

module bullet(input XVel, YVel,
					output XPos, YPos);
					
					
					