module bullet ( input Reset, frame_clk, //Faster clock needed
						input bullet_active,input angle,
                output [9:0]  BallX, BallY, BallS );
endmodule
					 
					 
